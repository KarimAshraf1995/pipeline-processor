library ieee;
use ieee.std_logic_1164.all;


entity Mux4 is 
	generic (width : integer := 16 );  
	port (S : in std_logic_vector(1 downto 0);
		A : in std_logic_vector (width-1 downto 0);
		B : in std_logic_vector (width-1 downto 0);
		C : in std_logic_vector (width-1 downto 0);
		D : in std_logic_vector (width-1 downto 0);
		F : out std_logic_vector(width-1 downto 0)
		);
end entity Mux4;


Architecture Mux4_Implementation of Mux4 is  
Begin 
	F <=  A when S="00" else
        B when S="01" else
        C when S="10"	else
        D;
  
end Architecture;
